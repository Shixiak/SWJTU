library verilog;
use verilog.vl_types.all;
entity Computer_vlg_vec_tst is
end Computer_vlg_vec_tst;
